//signed adder.
// passing two structures and one return str
module adder(a,b,c);
	input a,b;
	output c;
	// write the logic to add/subtract
	// WORK:
	// 1. see sign bits of a and b
	// 2. decide how to subtract
	// 3. put correct sign bit in c.
